LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;


PACKAGE definitions IS


---- globals
CONSTANT BUS_WIDTH : NATURAL := 32;
CONSTANT INST_WIDTH : NATURAL := 32;
CONSTANT ZEROS	: STD_LOGIC_VECTOR(31 downto 0) :=  "00000000000000000000000000000000";	
CONSTANT ONES	: STD_LOGIC_VECTOR(31 downto 0) :=  "11111111111111111111111111111111";	
CONSTANT ONES_MINUS	: STD_LOGIC_VECTOR(30 downto 0) :=  "1111111111111111111111111111111";	
CONSTANT ZEROS_MINUS	: STD_LOGIC_VECTOR(30 downto 0) :=  "0000000000000000000000000000000";	
CONSTANT ZEROS32	: STD_LOGIC_VECTOR(31 downto 0) :=  "00000000000000000000000000000000";		
	
	-- globals
--CONSTANT BUS_WIDTH : NATURAL := 8;
--CONSTANT INST_WIDTH : NATURAL := 32;
--CONSTANT ZEROS	: STD_LOGIC_VECTOR(7 downto 0) :=  "00000000";	
--CONSTANT ONES	: STD_LOGIC_VECTOR(7 downto 0) :=  "11111111";	
--CONSTANT ONES_MINUS	: STD_LOGIC_VECTOR(6 downto 0) :=  "1111111";	
--CONSTANT ZEROS_MINUS	: STD_LOGIC_VECTOR(6 downto 0) :=  "0000000";	
--CONSTANT ZEROS32	: STD_LOGIC_VECTOR(31 downto 0) :=  "00000000000000000000000000000000";	
END definitions;
